package lx32_all_pkg;
  import lx32_pkg::*;
  import branches_pkg::*;
endpackage

